netcdf test_hofx_sic_writer_out {
dimensions:
	N_QCF = 2 ;
	STRINGGRID = 1 ;
	STRINGJULD = 14 ;
	STRINGNAM = 8 ;
	STRINGTYP = 4 ;
	STRINGWMO = 8 ;
	N_OBS = 11 ;
	N_LEVELS = 1 ;
	N_VARS = 1 ;
	N_ENTRIES = 1 ;
	N_EXTRA = 1 ;
variables:
	char JULD_REFERENCE(STRINGJULD) ;
		JULD_REFERENCE:long_name = "Date of reference for julian days" ;
		JULD_REFERENCE:Conventions = "YYYYMMDDHHMMSS" ;
	char VARIABLES(N_VARS, STRINGNAM) ;
		VARIABLES:long_name = "List of variables in feedback files" ;
	char EXTRA(N_EXTRA, STRINGNAM) ;
	char ENTRIES(N_ENTRIES, STRINGNAM) ;
		ENTRIES:long_name = "List of additional entries for each variable in feedback files" ;
	double LATITUDE(N_OBS) ;
		LATITUDE:units = "degrees_north" ;
		LATITUDE:long_name = "latitude" ;
	double LONGITUDE(N_OBS) ;
		LONGITUDE:units = "degrees_east" ;
		LONGITUDE:long_name = "longitude" ;
	double DEPTH(N_OBS, N_LEVELS) ;
		DEPTH:units = "metre" ;
		DEPTH:long_name = "Depth" ;
	double JULD(N_OBS) ;
		JULD:units = "days since JULD_REFERENCE" ;
		JULD:long_name = "Julian day" ;
	char STATION_IDENTIFIER(N_OBS, STRINGWMO) ;
		STATION_IDENTIFIER:long_name = "Station identifier" ;
	char STATION_TYPE(N_OBS, STRINGTYP) ;
		STATION_TYPE:long_name = "Code instrument type" ;
	int DEPTH_QC(N_OBS, N_LEVELS) ;
		DEPTH_QC:long_name = "Quality on depth" ;
		DEPTH_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int DEPTH_QC_FLAGS(N_OBS, N_LEVELS, N_QCF) ;
		DEPTH_QC_FLAGS:long_name = "Quality on depth" ;
		DEPTH_QC_FLAGS:Conventions = "JEDI UFO QC flag conventions" ;
	int OBSERVATION_QC(N_OBS) ;
		OBSERVATION_QC:long_name = "Quality on observation" ;
		OBSERVATION_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int OBSERVATION_QC_FLAGS(N_OBS, N_QCF) ;
		OBSERVATION_QC_FLAGS:long_name = "Quality on observation" ;
		OBSERVATION_QC_FLAGS:Conventions = "JEDI UFO QC flag conventions" ;
	int POSITION_QC(N_OBS) ;
		POSITION_QC:long_name = "Quality on position" ;
		POSITION_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int POSITION_QC_FLAGS(N_OBS, N_QCF) ;
		POSITION_QC_FLAGS:long_name = "Quality on position" ;
		POSITION_QC_FLAGS:Conventions = "JEDI UFO QC flag conventions" ;
	int JULD_QC(N_OBS) ;
		JULD_QC:long_name = "Quality on date and time" ;
		JULD_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int JULD_QC_FLAGS(N_OBS, N_QCF) ;
		JULD_QC_FLAGS:long_name = "Quality on date and time" ;
		JULD_QC_FLAGS:Conventions = "JEDI UFO QC flag conventions" ;
	int ORIGINAL_FILE_INDEX(N_OBS) ;
		ORIGINAL_FILE_INDEX:long_name = "Index in original data file" ;
	double ICECONC_OBS(N_OBS, N_LEVELS) ;
		ICECONC_OBS:long_name = "ice area fraction" ;
		ICECONC_OBS:units = "Fraction" ;
		ICECONC_OBS:_FillValue = 99999. ;
	double ICECONC_Hx(N_OBS, N_LEVELS) ;
		ICECONC_Hx:long_name = "ice area fraction Hx" ;
		ICECONC_Hx:units = "Fraction" ;
		ICECONC_Hx:_FillValue = 99999. ;
	int ICECONC_QC_FLAGS(N_OBS, N_QCF) ;
		ICECONC_QC_FLAGS:_FillValue = 0 ;
		ICECONC_QC_FLAGS:long_name = "quality flags on ice area fraction" ;
		ICECONC_QC_FLAGS:Conventions = "OPS flag conventions" ;
	int ICECONC_LEVEL_QC_FLAGS(N_OBS, N_LEVELS, N_QCF) ;
		ICECONC_LEVEL_QC_FLAGS:_FillValue = 0 ;
		ICECONC_LEVEL_QC_FLAGS:long_name = "quality flags for each level on ice area fraction" ;
		ICECONC_LEVEL_QC_FLAGS:Conventions = "OPS flag conventions" ;
	int ICECONC_QC(N_OBS) ;
		ICECONC_QC:long_name = "quality on ice area fraction" ;
		ICECONC_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int ICECONC_LEVEL_QC(N_OBS, N_LEVELS) ;
		ICECONC_LEVEL_QC:_FillValue = 0 ;
		ICECONC_LEVEL_QC:long_name = "quality for each level on ice area fraction" ;
		ICECONC_LEVEL_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int ICECONC_IOBSI(N_OBS) ;
		ICECONC_IOBSI:long_name = "ORCA grid search I coordinate" ;
	int ICECONC_IOBSJ(N_OBS) ;
		ICECONC_IOBSJ:long_name = "ORCA grid search J coordinate" ;
	int ICECONC_IOBSK(N_OBS, N_LEVELS) ;
		ICECONC_IOBSK:long_name = "ORCA grid search K coordinate" ;
	char ICECONC_GRID(STRINGGRID) ;
		ICECONC_GRID:long_name = "ORCA grid search grid (T,U,V)" ;
	double MDT(N_OBS, N_LEVELS) ;
		MDT:long_name = "fake MDT" ;
		MDT:units = "fake metres" ;

// global attributes:
		:title = "NEMO observation operator output" ;
		:Convention = "NEMO unified observation operator output" ;
data:

 JULD_REFERENCE = "20210630120000" ;

 VARIABLES =
  "ICECONC " ;

 EXTRA =
  "MDT     " ;

 ENTRIES =
  "Hx      " ;

 LATITUDE = 82.029388, 62.43589, -65.285362, -51.879791, 41.894199, 
    22.651899, 3.3262999, -15.916, -35.2416, -54.483898, -73.726196 ;

 LONGITUDE = 168.338, 31.214951, -24.91501, -154.48199, 38.443001, -148.293, 
    25.115, -161.621, 11.787, -174.94901, -1.6849999 ;

 DEPTH =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 JULD = -1, -1, -1, -1, -0.5, -0.5, -0.5, -0.5, -0.5, -0.5, -0.5 ;

 STATION_IDENTIFIER =
  "        ",
  "        ",
  "        ",
  "        ",
  "        ",
  "        ",
  "        ",
  "        ",
  "        ",
  "        ",
  "        " ;

 STATION_TYPE =
  "0   ",
  "0   ",
  "0   ",
  "0   ",
  "0   ",
  "0   ",
  "0   ",
  "0   ",
  "0   ",
  "0   ",
  "0   " ;

 DEPTH_QC =
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _ ;

 DEPTH_QC_FLAGS =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

 OBSERVATION_QC = 4, 4, 4, 1, 4, 1, 4, 1, 1, 1, 4 ;

 OBSERVATION_QC_FLAGS =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

 POSITION_QC = _, _, _, _, _, _, _, _, _, _, _ ;

 POSITION_QC_FLAGS =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

 JULD_QC = _, _, _, _, _, _, _, _, _, _, _ ;

 JULD_QC_FLAGS =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

 ORIGINAL_FILE_INDEX = _, _, _, _, _, _, _, _, _, _, _ ;

 ICECONC_OBS =
  0,
  _,
  0.99629998,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 ICECONC_Hx =
  0.495,
  _,
  0,
  0,
  _,
  0,
  _,
  0,
  0,
  0,
  _ ;

 ICECONC_QC_FLAGS =
  68, _,
  1, _,
  68, _,
  64, _,
  1, _,
  64, _,
  1, _,
  64, _,
  64, _,
  64, _,
  1, _ ;

 ICECONC_LEVEL_QC_FLAGS =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

 ICECONC_QC = 4, 4, 4, 1, 4, 1, 4, 1, 1, 1, 4 ;

 ICECONC_LEVEL_QC =
  4,
  4,
  4,
  1,
  4,
  1,
  4,
  1,
  1,
  1,
  4 ;

 ICECONC_IOBSI = _, _, _, _, _, _, _, _, _, _, _ ;

 ICECONC_IOBSJ = _, _, _, _, _, _, _, _, _, _, _ ;

 ICECONC_IOBSK =
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _ ;

 ICECONC_GRID = "T" ;

 MDT =
  0,
  99999,
  0.99629998,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;
}
