netcdf test_hofx_profiles_writer_out {
dimensions:
	N_QCF = 2 ;
	STRINGGRID = 1 ;
	STRINGJULD = 14 ;
	STRINGNAM = 8 ;
	STRINGTYP = 4 ;
	STRINGWMO = 8 ;
	N_OBS = 1 ;
	N_LEVELS = 10 ;
	N_VARS = 1 ;
	N_ENTRIES = 1 ;
variables:
	char JULD_REFERENCE(STRINGJULD) ;
		JULD_REFERENCE:long_name = "Date of reference for julian days" ;
		JULD_REFERENCE:Conventions = "YYYYMMDDHHMMSS" ;
	char VARIABLES(N_VARS, STRINGNAM) ;
		VARIABLES:long_name = "List of variables in feedback files" ;
	char ENTRIES(N_ENTRIES, STRINGNAM) ;
		ENTRIES:long_name = "List of additional entries for each variable in feedback files" ;
	double LATITUDE(N_OBS) ;
		LATITUDE:units = "degrees_north" ;
		LATITUDE:long_name = "latitude" ;
	double LONGITUDE(N_OBS) ;
		LONGITUDE:units = "degrees_east" ;
		LONGITUDE:long_name = "longitude" ;
	double DEPTH(N_OBS, N_LEVELS) ;
		DEPTH:units = "metre" ;
		DEPTH:long_name = "Depth" ;
	double JULD(N_OBS) ;
		JULD:units = "days since JULD_REFERENCE" ;
		JULD:long_name = "Julian day" ;
	char STATION_IDENTIFIER(N_OBS, STRINGWMO) ;
		STATION_IDENTIFIER:long_name = "Station identifier" ;
	char STATION_TYPE(N_OBS, STRINGTYP) ;
		STATION_TYPE:long_name = "Code instrument type" ;
	int DEPTH_QC(N_OBS, N_LEVELS) ;
		DEPTH_QC:long_name = "Quality on depth" ;
		DEPTH_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int DEPTH_QC_FLAGS(N_OBS, N_LEVELS, N_QCF) ;
		DEPTH_QC_FLAGS:long_name = "Quality on depth" ;
		DEPTH_QC_FLAGS:Conventions = "OPS flag conventions" ;
	int OBSERVATION_QC(N_OBS) ;
		OBSERVATION_QC:long_name = "Quality on observation" ;
		OBSERVATION_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int OBSERVATION_QC_FLAGS(N_OBS, N_QCF) ;
		OBSERVATION_QC_FLAGS:long_name = "Quality on observation" ;
		OBSERVATION_QC_FLAGS:Conventions = "OPS flag conventions" ;
	int POSITION_QC(N_OBS) ;
		POSITION_QC:long_name = "Quality on position" ;
		POSITION_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int POSITION_QC_FLAGS(N_OBS, N_QCF) ;
		POSITION_QC_FLAGS:long_name = "Quality on position" ;
		POSITION_QC_FLAGS:Conventions = "OPS flag conventions" ;
	int JULD_QC(N_OBS) ;
		JULD_QC:long_name = "Quality on date and time" ;
		JULD_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int JULD_QC_FLAGS(N_OBS, N_QCF) ;
		JULD_QC_FLAGS:long_name = "Quality on date and time" ;
		JULD_QC_FLAGS:Conventions = "OPS flag conventions" ;
	int ORIGINAL_FILE_INDEX(N_OBS) ;
		ORIGINAL_FILE_INDEX:long_name = "Index in original data file" ;
	double POTM_OBS(N_OBS, N_LEVELS) ;
		POTM_OBS:long_name = "sea water potential temperature" ;
		POTM_OBS:units = "degrees Celsius" ;
		POTM_OBS:_FillValue = 99999. ;
	double POTM_Hx(N_OBS, N_LEVELS) ;
		POTM_Hx:long_name = "sea water potential temperature Hx" ;
		POTM_Hx:units = "degrees Celsius" ;
		POTM_Hx:_FillValue = 99999. ;
	int POTM_QC_FLAGS(N_OBS, N_QCF) ;
		POTM_QC_FLAGS:_FillValue = 0 ;
		POTM_QC_FLAGS:long_name = "quality flags on sea water potential temperature" ;
		POTM_QC_FLAGS:Conventions = "OPS flag conventions" ;
	int POTM_LEVEL_QC_FLAGS(N_OBS, N_LEVELS, N_QCF) ;
		POTM_LEVEL_QC_FLAGS:_FillValue = 0 ;
		POTM_LEVEL_QC_FLAGS:long_name = "quality flags for each level on sea water potential temperature" ;
		POTM_LEVEL_QC_FLAGS:Conventions = "OPS flag conventions" ;
	int POTM_QC(N_OBS) ;
		POTM_QC:long_name = "quality on sea water potential temperature" ;
		POTM_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int POTM_LEVEL_QC(N_OBS, N_LEVELS) ;
		POTM_LEVEL_QC:_FillValue = 0 ;
		POTM_LEVEL_QC:long_name = "quality for each level on sea water potential temperature" ;
		POTM_LEVEL_QC:Conventions = "U.S. Integrated Ocean Observing System, 2017. Manual for the Use of Real-Time Oceanographic Data Quality Control Flags, Version 1.1" ;
	int POTM_IOBSI(N_OBS) ;
		POTM_IOBSI:long_name = "ORCA grid search I coordinate" ;
	int POTM_IOBSJ(N_OBS) ;
		POTM_IOBSJ:long_name = "ORCA grid search J coordinate" ;
	int POTM_IOBSK(N_OBS, N_LEVELS) ;
		POTM_IOBSK:long_name = "ORCA grid search K coordinate" ;
	char POTM_GRID(STRINGGRID) ;
		POTM_GRID:long_name = "ORCA grid search grid (T,U,V)" ;

// global attributes:
		:title = "NEMO observation operator output" ;
		:Convention = "NEMO unified observation operator output" ;
data:

 JULD_REFERENCE = "19500101000000" ;

 VARIABLES =
  "POTM    " ;

 ENTRIES =
  "Hx      " ;

 LATITUDE = 35 ;

 LONGITUDE = -40 ;

 DEPTH =
  0, 1, 2, 3, 4, 5, 10, 100, 200, 1000 ;

 JULD = 26113.5 ;

 STATION_IDENTIFIER =
  "20190615" ;

 STATION_TYPE =
  "    " ;

 DEPTH_QC =
  _, _, _, _, _, _, _, _, _, _ ;

 DEPTH_QC_FLAGS =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

 OBSERVATION_QC = 0 ;

 OBSERVATION_QC_FLAGS =
  _, _ ;

 POSITION_QC = _ ;

 POSITION_QC_FLAGS =
  _, _ ;

 JULD_QC = _ ;

 JULD_QC_FLAGS =
  _, _ ;

 ORIGINAL_FILE_INDEX = _ ;

 POTM_OBS =
  12.3000001907349, 12.3999996185303, 12.8999996185303, _, 11.6999998092651, 
    10.3000001907349, 10.6999998092651, 9.30000019073486, 9.10000038146973, _ ;

 POTM_Hx =
  18.1944444613818, 12.3999996185303, 12.8999996185303, _, 11.6999998092651, 
    10.3000001907349, 10.6999998092651, 9.30000019073486, 9.10000038146973, _ ;

 POTM_QC_FLAGS =
  _, _ ;

 POTM_LEVEL_QC_FLAGS =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;

 POTM_QC = 1 ;

 POTM_LEVEL_QC =
  1, 1, 4, 4, 1, 4, 1, 1, 4, 4 ;

 POTM_IOBSI = _ ;

 POTM_IOBSJ = _ ;

 POTM_IOBSK =
  _, _, _, _, _, _, _, _, _, _ ;

 POTM_GRID = "T" ;
}
